entity test is
port();
end entity
