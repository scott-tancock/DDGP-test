entity test is
port(
	clk : in std_logic;
	rst : in std_logic);
end entity
