entity tb_test is
port();
end entity;
